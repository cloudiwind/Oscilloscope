`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: NUS ECE
// Engineer: Shahzor Ahmad
// 
// Create Date: 02.10.2015 14:31:19
// Design Name: 
// Module Name: SCOPE_TOP
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////////


module SCOPE_TOP(

    input CLK,                  // main system clock, 100MHz
        
    input btnL,                 // buttons
    input btnR,
    input btnU,
    input btnC,
    input btnD,    

    input ADC_IN_P,             // differential +ve & -ve analog inputs to ADC
    input ADC_IN_N,  
    
    input TRIGGER,              // toggle triggering
    input TRIGGER_TYPE,        // changing wave types (square, sin, tri)
    
    output reg[3:0] VGA_RED,    // RGB outputs to VGA connector (4 bits per channel gives 4096 possible colors)
    output reg[3:0] VGA_GREEN,
    output reg[3:0] VGA_BLUE,
    output reg VGA_VS,          // horizontal & vertical sync outputs to VGA connector
    output reg VGA_HS,
    
    output [11:0] led           // debug LEDs    
    
    );   
         
    //-------------------------------------------------------------------------
    
    wire CLK_MAIN = CLK ;   // this is just a renaming (simply a short-circuit, or two names for the same trace/route)           
       
        
    //-------------------------------------------------------------------------
    
    //         INSTANTITATE EXTERNAL MODULES FOR VGA CONTROL
    
    // Note the VGA controller is configured to produce a 1024 x 1280 pixel resolution
    //-------------------------------------------------------------------------
    
    // PIXEL CLOCK GENERATOR 
    wire CLK_VGA ;          // pixel/VGA clock is generated by MMCM/PLL via external VHDL code (108MHz)    
    clk_wiz_0 PIXEL_CLOCK_GENERATOR( 
            CLK_MAIN,   // 100 MHz
            CLK_VGA     // 108 MHz
        ) ;     
    
    
    // VGA SIGNALS (as output by VGA controller (vga_ctrl.vhd))
    wire VGA_horzSync ;
    wire VGA_vertSync ;
    wire VGA_active ;
    wire[11:0] VGA_horzCoord ;
    wire[11:0] VGA_vertCoord ;
        // it is not required but good practice to declare single-bit wires
        // it is required to declare multi-bit wires (bus) before use    
    
    // VGA CONTROLLER    
    vga_ctrl VGA_CONTROLLER(
            CLK_VGA,
            VGA_horzSync,
            VGA_vertSync,
            VGA_active,  
            VGA_horzCoord,  
            VGA_vertCoord  
        ) ; 
        // - VGA_horzCoord changes at a rate of 108 MHz (CLK_VGA) to traverse each pixel in a row, while VGA_vertCoord changes at a rate of ~63.98 KHz to 
        // scan each row one by one and back to the top. These tech details are handled by vga_ctrl.vhd. One only needs to make use of these coordinates 
        // to output whatever they want at desired pixel locations. 
        // 
        // - VGA_active is a binary indicator specifying when VGA_horzCoord, VGA_vertCoord are valid (i.e., with the 1024 x 1280 pixel screen). For technical 
        // reasons the said coordinates do go outside this screen area for a short while and no VGA signal should be output during this time (it will and does
        // mess up the display). 
        //
        // - hence, VGA_active, VGA_horzCoord and VGA_vertCoord may be used in conjunction with each other to generate VGA_RED, VGA_GREEN, VGA_BLUE. The Sync
        // signals should be output to the VGA port as well, and are responsible to generate the raster scan on the screen       


    //-------------------------------------------------------------------------
                                    
    //                      SAMPLING VIA ADC 
    
    // On-chip ADC is clocked at [ inv(inv(CLK_ADC/4)*26) = 961.538 KHZ ], 
    // where CLK_ADC is the clock passed to ADC (in this case CLK_ADC = CLK_MAIN = 100MHz)
    
    // The on-chip ADC is 12-bit. We employ the most significant 8 bits to keep things simple
    
    //-------------------------------------------------------------------------
    
    wire [7:0] ADC_SAMPLE ; // the latest value as sampled via ADC
    ADC_sampler SAMPLER(CLK_MAIN, ADC_IN_P, ADC_IN_N, ADC_SAMPLE ) ; // sampling at 961.538 KHZ
        // Either lines # 104-105 OR lines # 129-136 should be used at a time

    //assign led[7:0] = ADC_SAMPLE ; 
        // the sampled 8-bit value reflects on 8 LEDs. Every time ADC_SAMPLE changes 
        // (and that happens at 961.538KHz!), this assignment is triggered again 
      
    
    //-------------------------------------------------------------------------
                                        
    //                  SIMULATE SAMPLING VIA ADC 
    
    // In the absence of a signal generator (e.g., when working at home), you may use 
    // the following code instead of the above, i.e., COMMENT out lines # 104-105, 
    // UN-COMMENT lines # 129-136
    
    // A square wave at 1Hz is generated via a clock-divider module, and serves as our 
    // 'analog' signal to be sampled.
    //-------------------------------------------------------------------------
    
    wire CLK_SYNTH_SQUARE ; 
    clock_divider GEN_CLK_SYNTH_SQUARE( CLK_MAIN, 1'b0, 28'H2FAF080, CLK_SYNTH_SQUARE ) ; 
        // Synthesize a 1Hz waveform given 100MHz clock          
/*
    reg [7:0] ADC_SAMPLE ; // the latest value as sampled via ADC
    always@(posedge CLK_MAIN) // sample the synthesized waveform at 100 MHz
        begin
            if( CLK_SYNTH_SQUARE )
                ADC_SAMPLE <= 255 ;
            else
                ADC_SAMPLE <= 0 ;        
        end       
*/
     // this LED blinks at 1 Hz (just for visualization)
     reg LED_DEBUG = 0 ;
        // signals on LHS of assignments in 'always' blocks must be declared as reg before use
//     always@(posedge CLK_SYNTH_SQUARE)
//        begin
//            LED_DEBUG <= !LED_DEBUG ;
//        end
//     assign led[8] = LED_DEBUG ; 
     
//     clock_divider GEN_CLK_SYNTH_TRI(CLK_MAIN, 1'b0, 28'H004F080, CLK2);
     
//     reg dirn = 0;
//     reg [7:0] ADC_SAMPLE = 0;
     
//     always @ (posedge CLK2) begin
//        if (!dirn)
//            ADC_SAMPLE = ADC_SAMPLE + 1;
//        else
//            ADC_SAMPLE = ADC_SAMPLE - 1;
//        if (ADC_SAMPLE == 8'b11111111 || ADC_SAMPLE == 0)
//            dirn = ~dirn;
//     end   
               
    //-------------------------------------------------------------------------
                                    
    //        SELECTING SAMPLING FREQUENCY (ESSENTIALLY, TIME/DIV)
    
    // this configures the CLK_SUBSAMPLE (fs)
    
    // NOTE: currently CLK_SUBSAMPLE_ID has been hard-coded to 0, and no provision
    // is made to modify it at FPGA run-time
    //-------------------------------------------------------------------------
    
    reg [2:0] CLK_SUBSAMPLE_ID = 0 ; 
        
    reg [27:0] LOAD_VALUE_SUBSAMPLE ;
        // we generate CLK_SUBSAMPLE from CLK_MAIN 
    
    always@(posedge CLK_MAIN)
        case(CLK_SUBSAMPLE_ID)
            0:  LOAD_VALUE_SUBSAMPLE <= 28'd500000 ;    // CLK_SUBSAMPLE = 100 Hz => TIME/DIV = 0.8 sec/div
            1:  LOAD_VALUE_SUBSAMPLE <= 28'd125000 ;    // CLK_SUBSAMPLE = 400 Hz => TIME/DIV = 0.2 sec/div 
            2:  LOAD_VALUE_SUBSAMPLE <= 28'd62500 ;     // CLK_SUBSAMPLE = 800 Hz => TIME/DIV = 0.1 sec/div
            3:  LOAD_VALUE_SUBSAMPLE <= 28'd50000 ;     // CLK_SUBSAMPLE = 1 KHz => TIME/DIV = 
            4:  LOAD_VALUE_SUBSAMPLE <= 28'd31250 ;     // CLK_SUBSAMPLE = 1600 Hz => TIME/DIV = 50 ms/div 
            5:  LOAD_VALUE_SUBSAMPLE <= 28'd6250 ;      // CLK_SUBSAMPLE = 8 KHz => TIME/DIV = 10 ms/div 
            6:  LOAD_VALUE_SUBSAMPLE <= 28'd625 ;       // CLK_SUBSAMPLE = 80 KHz => TIME/DIV = 1 ms/div      
            7:  LOAD_VALUE_SUBSAMPLE <= 28'd62 ;        // CLK_SUBSAMPLE = 806.451 KHz => TIME/DIV = 0.0992 ms/div 
        endcase
            // Each LOAD_VALUE_SUBSAMPLE defines the stated CLK_SUBSAMPLE (sampling frequency fs). 
            // The TIME/DIV values, however, assume the 1280 horizontal pixels on the screen are divided into 16 equal DIVISIONS of 80 px each 
                      
    
    wire CLK_SUBSAMPLE, CLK_2 ;    // sub-sampling rate for ADC output samples
                            // It essentially defines time/div 
                            
                            // Use CLK_SUBSAMPLE to clock your bank of shift registers below
                            // Use CLK_SUBSAMPLE to clock your trigger process if you implement one   
                            
                            // For all practical purposes, this can be taken to be our fs (sampling frequency) as described in the manual
                            // We could have modified ADC sampling frequency, but give the long formula to dervie it from CLK_MAIN (see line 96),
                            // we're better off sub-sampling to achieve flexible sampling frequencies and corresponding time/div configurations
                                                        
                                                     
    clock_divider GEN_CLK_SUBSAMPLE( CLK_MAIN, 1'b0, LOAD_VALUE_SUBSAMPLE, CLK_SUBSAMPLE ) ;
    clock_divider GEN_CLK_2( CLK_MAIN, 1'b0, 28'd4000000, CLK_2 ) ;
//    clock_divider GEN_CLK_CURSOR (CLK_MAIN, 1'b0, 28'd50, CLK_CURSOR);

        // note as many times you instantiate a module in HDL, that many times it will replicate the actual hardware on the FPGA 
        // so there are two physical clock_divider circuits in our design    
    
    switch_debouncer TRIG_DEBOUNCER( CLK_MAIN, TRIGGER, TRIGGER_DB ) ;
    switch_debouncer TRIG_TYPE_DEBOUNCER (CLK_MAIN, TRIGGER_TYPE, TRIGGER_TYPE_DB); 
    
    button_debouncer DEBOUNCE_LHS (CLK_2, btnL, LHS_DEBOUNCE); 
    button_debouncer DEBOUNCE_RHS (CLK_2, btnR, RHS_DEBOUNCE); 
    button_debouncer DEBOUNCE_TOP (CLK_2, btnU, TOP_DEBOUNCE); 
    button_debouncer DEBOUNCE_BTM (CLK_2, btnC, BTM_DEBOUNCE); 
        
        // you may implement debounce in switch_debouncer.vhd as an extension feature
    CHANGE_SPEED showSpeed(CLK_SUBSAMPLE_ID, OP0, OP1, OP2, OP3, OP4, OP5, OP6, OP7);
    
    wire [1:0] ctrl ; 
//    FSM_inc_dec FSM1( CLK_MAIN, btnL, btnR, ctrl ) ;        // use if you don't implement debounce, but would like to write an FSM
    //assign led[13:12] = ctrl;
    FSM_inc_dec FSM1(CLK_2, TOP_DEBOUNCE, BTM_DEBOUNCE, ctrl) ;  // use if you've implemented debounce, and now would also like to implement FSM
    
    always @(posedge CLK_2) begin
        if( ctrl == 2'b01 && CLK_SUBSAMPLE_ID < 7 )
            CLK_SUBSAMPLE_ID <= CLK_SUBSAMPLE_ID + 1 ;
        else if (ctrl == 2'b10 && CLK_SUBSAMPLE_ID > 0)
            CLK_SUBSAMPLE_ID <= CLK_SUBSAMPLE_ID - 1 ;
    end        
        // you may implement a FSM in FSM_inc_dec.vhd as an extension feature
        // This FSM should output a 2-bit control sisgnal
        //      00 -- do nothing
        //      01 -- increment CLK_SUBSAMPLE_ID
        //      10 -- decrement CLK_SUBSAMPLE_ID

    //assign ctrl = 0 ; // remove this if you implement your FSM

    // this process increments / decrements CLK_SUBSAMPLE_ID depending on ctrl        
//    always@(posedge CLK_MAIN)
//        begin
//            if( ctrl == 2'b01 )
//                CLK_SUBSAMPLE_ID = CLK_SUBSAMPLE_ID + 1 ;
//            else if (ctrl == 2'b10)
//                CLK_SUBSAMPLE_ID = CLK_SUBSAMPLE_ID - 1 ;
//        end
     

    assign led[11:9] = CLK_SUBSAMPLE_ID ;  
        // leds[11:9] provide a visual indication of CLK_SUBSAMPLE_ID at all times    
  
    
    //-------------------------------------------------------------------------
                                    
    //               UPDATE DISPLAY_MEM @ CLK_SUBSAMPLE
    
    // DISPLAY_MEM is a bank of 1280 shift registers
    
    // shift all samples one position to the left in memory, and  
    // store the latest ADC sample in the right/left most position    
    //-------------------------------------------------------------------------

    reg [7:0] DISPLAY_MEM[0:1279] ;
    //reg [7:0] DISPLAY_NEW[0:1279] ; 
    reg [7:0] DISPLAY_TEMP[0:1279] ;
        // display memory - store samples here and output them on screen
        
    // TOOD:    implement Verilog here that treats DISPLAY_MEM as a bank of 
    //          1280 shift registers, each 8-bit wide. The latest sample should 
    //          be stored in the right (or left)-most register, while contents of
    //          all the other registers should be shifted to the neighboring register
    //          on the right (respectively, left). 
    //          
    //          This process of bringing in a new sample from the right/left while 
    //          shifting all the other samples should be done in a single clock cycle 
    //          (use CLK_SUBSAMPLE)

    integer i;
    integer j;
    
    // Coupled with start-stop function
    always @ (posedge CLK_SUBSAMPLE) begin
       if (~btnD) begin
           for( i = 0; i<1279 ; i = i+1 ) begin
                    DISPLAY_TEMP[i+1] <= DISPLAY_TEMP[i];
           end
           DISPLAY_TEMP[0] <= ADC_SAMPLE;
        end 
    end


    // TRIGGER_TYPE_DB toggles between square waves and non-square waves
    always @ (posedge CLK_SUBSAMPLE) begin
            if ((ADC_SAMPLE >= 20 && ADC_SAMPLE > DISPLAY_TEMP[1] && TRIGGER_DB && TRIGGER_TYPE_DB) ||
            (ADC_SAMPLE == 20 && ADC_SAMPLE > DISPLAY_TEMP[1] && TRIGGER_DB && ~TRIGGER_TYPE_DB) || ~TRIGGER_DB ) begin
            
                for( j = 0; j<1280 ; j = j+1 ) begin
                    DISPLAY_MEM[j] <= DISPLAY_TEMP[j];
                end
            end
        end    
   
    
    
    
    //-------------------------------------------------------------------------
                
    //                  DRAWING WAVEFORM ON SCREEN
    
    // waveform is drawn using its samples from display memory
    //-------------------------------------------------------------------------       
           
    wire[3:0] VGA_GREEN_WAVEFORM =                         //Original 511+128
                ((VGA_horzCoord < 1280) & (VGA_vertCoord == ((511+128) - DISPLAY_MEM[VGA_horzCoord]))) //||
//                ((VGA_horzCoord < 1280) & (VGA_vertCoord == ((511+128) - DISPLAY_NEW[VGA_horzCoord])))
                    ? 4'hF : 0 ;             
                
    //-------------------------------------------------------------------------
        
    //                  DRAWING GRID LINES ON SCREEN
    
    // Grid lines are drawn at pixels # 320, 640, 960 along the x-axis, and
    // pixels # 256, 512, 768 along the y-axis
    
    // Note the VGA controller is configured to produce a 1024 x 1280 pixel resolution
    //-------------------------------------------------------------------------
    
    wire CONDITION_FOR_GRID = (VGA_horzCoord%80 == 79) || (VGA_vertCoord%64 == 63);        
           
    wire CONDITION_FOR_TICKS = ((VGA_horzCoord%16 == 15) && (509 <= VGA_vertCoord && VGA_vertCoord <= 513)) ||
                               ((VGA_vertCoord%8 == 7) && (637 <= VGA_horzCoord && VGA_horzCoord <= 641)); 
          
    //wire CONDITION_FOR_GRID = (VGA_horzCoord == 319) || (VGA_horzCoord == 639) || (VGA_horzCoord == 959) ||
    //                (VGA_vertCoord == 255) || (VGA_vertCoord == 511) || (VGA_vertCoord == 767) ;
    
    wire[3:0] VGA_RED_GRID = (CONDITION_FOR_GRID || CONDITION_FOR_TICKS) ? 0 : 4'h7 ;
    wire[3:0] VGA_GREEN_GRID = (CONDITION_FOR_GRID || CONDITION_FOR_TICKS) ? 0 : 4'h3 ;
    wire[3:0] VGA_BLUE_GRID = (CONDITION_FOR_GRID || CONDITION_FOR_TICKS) ? 0 : 4'h5 ;
        // if true, a black pixel is put at coordinates (VGA_horzCoord, VGA_vertCoord), 
        // else a cyan background is generated, characteristic of oscilloscopes! 
        
    // TOOD:    Draw grid lines at every 80-th pixel along the horizontal axis, and every 64th pixel
    //          along the vertical axis. This gives us a 16x16 grid on screen. 
    //          
    //          Further draw ticks on the central x and y grid lines spaced 16 and 8 pixels apart in the 
    //          horizontal and vertical directions respectively. This gives us 5 sub-divisions per division 
    //          in the horizontal and 8 sub-divisions per divsion in the vertical direction   
    
    ConditionForMyName MY_NAME (VGA_vertCoord, VGA_horzCoord, CONDITION_FOR_MY_NAME);
    wire [3:0] VGA_FOR_MY_NAME = (CONDITION_FOR_MY_NAME) ? 4'hF : 0;
 
    ConditionFor0 ZERO (VGA_vertCoord, VGA_horzCoord, CDN_0);
    ConditionFor1 ONE (VGA_vertCoord, VGA_horzCoord, CDN_1);
    ConditionFor2 TWO (VGA_vertCoord, VGA_horzCoord, CDN_2);
    ConditionFor3 THREE (VGA_vertCoord, VGA_horzCoord, CDN_3);
    ConditionFor4 FOUR (VGA_vertCoord, VGA_horzCoord, CDN_4);
    ConditionFor5 FIVE (VGA_vertCoord, VGA_horzCoord, CDN_5);
    ConditionFor6 SIX (VGA_vertCoord, VGA_horzCoord, CDN_6);
    ConditionFor7 SEVEN (VGA_vertCoord, VGA_horzCoord, CDN_7);
    
    wire[3:0] VGA_0 = (CDN_0 & OP0) ? 4'hF : 0;
    wire[3:0] VGA_1 = (CDN_1 & OP1) ? 4'hF : 0;
    wire[3:0] VGA_2 = (CDN_2 & OP2) ? 4'hF : 0;
    wire[3:0] VGA_3 = (CDN_3 & OP3) ? 4'hF : 0;
    wire[3:0] VGA_4 = (CDN_4 & OP4) ? 4'hF : 0;
    wire[3:0] VGA_5 = (CDN_5 & OP5) ? 4'hF : 0;
    wire[3:0] VGA_6 = (CDN_6 & OP6) ? 4'hF : 0;
    wire[3:0] VGA_7 = (CDN_7 & OP7) ? 4'hF : 0;
 
    //-------------------------------------------------------------------------
    
    //              SYNCHRONOUS OUTPUT OF VGA SIGNALS
    
    //-------------------------------------------------------------------------
    
    // COMBINE ALL OUTPUTS ON EACH CHANNEL
    wire[3:0] VGA_RED_CHAN = VGA_RED_GRID ;
    wire[3:0] VGA_GREEN_CHAN = VGA_GREEN_GRID | VGA_GREEN_WAVEFORM | VGA_FOR_MY_NAME |
                               VGA_0 | VGA_1 | VGA_2 | VGA_3 | VGA_4 | VGA_5 | VGA_6 | VGA_7;; 
    wire[3:0] VGA_BLUE_CHAN = VGA_BLUE_GRID | VGA_FOR_MY_NAME |
                                VGA_0 | VGA_1 | VGA_2 | VGA_3 | VGA_4 | VGA_5 | VGA_6 | VGA_7;  


    // CLOCK THEM OUT
    always@(posedge CLK_VGA)
        begin      
        
            VGA_RED <= {VGA_active, VGA_active, VGA_active, VGA_active} & VGA_RED_CHAN ;  
            VGA_GREEN <= {VGA_active, VGA_active, VGA_active, VGA_active} & VGA_GREEN_CHAN ; 
            VGA_BLUE <= {VGA_active, VGA_active, VGA_active, VGA_active} & VGA_BLUE_CHAN ; 
                // VGA_active turns off output to screen if scan lines are outside the active screen area
            
            VGA_HS <= VGA_horzSync ;
            VGA_VS <= VGA_vertSync ;
            
        end
endmodule
